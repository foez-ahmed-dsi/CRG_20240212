//////////////////////////////////////////////////////////////////////////////////////////////////
// Name: Sadman Ishrak
// Email: sadmanishrak.work@gmail.com
//////////////////////////////////////////////////////////////////////////////////////////////////
module upper_module
(
    input logic pll_i [4],
    input logic [1:0] sel_i,
    input logic arst_ni,
    input logic en_i,
    output logic clk_out_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

    logic clk_mux_out_net;




//////////////////////////////////////////////////////////////////////////////////////////////////
// INSTANCES
//////////////////////////////////////////////////////////////////////////////////////////////////

    clk_mux_4x1 clk_mux_inst (
        .sel_i(sel_i),
        .pll_i(pll_i),
        .pll_o(clk_mux_out_net)
    );

    clk_gate clk_gate_inst (
        .en_i(en_i),
        .clk_i(clk_mux_out_net),
        .arst_ni(arst_ni),
        .pll_o(clk_out_o)
    );

endmodule
