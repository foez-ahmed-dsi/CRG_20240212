//////////////////////////////////////////////////////////////////////////////////////////////////
// Name: Sadman Ishrak
// Email: sadmanishrak.work@gmail.com
//////////////////////////////////////////////////////////////////////////////////////////////////
module upper_module
(
    input logic [3:0] pll_i,
    input logic [1:0] sel_i,
    input logic arst_n_i,
    input logic en_i,
    output logic clk_out_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

    logic clk_mux_out_net;




//////////////////////////////////////////////////////////////////////////////////////////////////
// INSTANCES
//////////////////////////////////////////////////////////////////////////////////////////////////

    clk_mux_4X1 clk_mux_inst (
        .sel_i(sel_i),
        .pll_i(pll_i),
        .pll_o(clk_mux_out_net)
    );

    clock_gate clk_gate_inst (
        .en_i(en_i),
        .clk_i(clk_mux_out_net),
        .arstn_i(arst_n_i),
        .pll_o(clk_out)
    );

endmodule
