//////////////////////////////////////////////////////////////////////////////////////////////////
// Name: Sadman Ishrak
// Email: sadmanishrak.work@gmail.com
//////////////////////////////////////////////////////////////////////////////////////////////////

module clk_mux_2x1(
    input logic sel_i,
    input logic pll_1_i,
    input logic pll_2_i,
    output logic clk_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

  logic q1, q2;


//////////////////////////////////////////////////////////////////////////////////////////////////
// SEQUENTIAL
//////////////////////////////////////////////////////////////////////////////////////////////////

  always @ (posedge pll_1_i) begin
    q1 <= ~sel_i && ~q2;
  end

  always @ (posedge pll_2_i) begin
    q2 <= sel_i && ~q1;
  end

//////////////////////////////////////////////////////////////////////////////////////////////////
// COMBINATIONAL
//////////////////////////////////////////////////////////////////////////////////////////////////

  assign clk_o = (q1 && pll_1_i) || (q2 && pll_2_i);

endmodule
