module rst_out
