// Description here
// ### Author : Nazmus Sakib (nazmus.sakib.punno@dsinnovators.com)

`include "clocking.svh"

module arst_no_tb;
  `define ENABLE_DUMPFILE

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-IMPORTS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // bring in the testbench essentials functions and macros
  `include "tb_ess.svh"

  //}}}


  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // generates static task start_clk_i with tHigh:4ns tLow:6ns
  `CREATE_CLK(ref_clk_i, 5ns, 5ns)
  logic glob_arst_ni=1;
  logic arst_req_i=0;
  logic arst_no;

  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////



  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////
  arst_no u_arst_no(
    .glob_arst_ni(glob_arst_ni),
    .arst_req_i(arst_req_i),
    .ref_clk_i(ref_clk_i),
    .arst_n(arst_n)
  );


  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////
 
  task static rand_arst_req_i(realtime unit_time = 1ns, int unsigned min = 50,
                          int unsigned max = 200);
    fork
      forever begin
        #(unit_time * $urandom_range(min, max));
        arst_req_i<= ($urandom_range(0,99)<15);
      end
    join_none
  endtask

  task static rand_glob_arst_ni(realtime unit_time = 1ns, int unsigned min = 50,
                          int unsigned max = 200);
    fork
      forever begin
        #(unit_time * $urandom_range(min, max));
        glob_arst_ni<= ($urandom_range(0,99)<95);
      end
    join_none
  endtask

  task static apply_reset();  //{{{
    #20ns;
    glob_arst_ni <= 0;
    #30ns;
    glob_arst_ni <= 1;
    #100ns;
  endtask  //}}}

  //}}}

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS{{{
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial{{{
    apply_reset();
    start_ref_clk_i();
    rand_arst_req_i();
    rand_glob_arst_ni();
    

    @(posedge clk_i);
    result_print(1, "This is a PASS");
    @(posedge clk_i);
    result_print(0, "And this is a FAIL");

    $finish;

  end  //}}}

  //}}}

endmodule
