//////////////////////////////////////////////////////////////////////////////////////////////////
// Name : Shahid Uddin Ahmed
// Email : shahid.ahmed@dsinnovators.com
//////////////////////////////////////////////////////////////////////////////////////////////////


module edge_detector(
    input logic e_data_i,
    input logic clk_ref_i,
    output logic edge_out_bar_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

    logic d_2, q_bar_1;

//////////////////////////////////////////////////////////////////////////////////////////////////
// SEQUENTIAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @ (posedge clk_ref_i) begin
        q_bar_1 <= ~(e_data_i);
    end

    always_ff @ (posedge clk_ref_i) begin
        edge_out_bar_o <= ~d_2;
    end

//////////////////////////////////////////////////////////////////////////////////////////////////
// COMBINATIONAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    always_comb begin
        d_2 = ~(q_bar_1 | e_data_i);
    end



endmodule

