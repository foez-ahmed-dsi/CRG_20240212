////////////////////////////////////////////////////////////////////////////////
//
//  Author - Sadman Ishrak
//  Email - sadmaishrak.work@gmail.com
//
////////////////////////////////////////////////////////////////////////////////
module clk_gate(
    input logic en_i,
    input logic clk_i,
    input logic arst_ni,
    output logic pll_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

    logic clk_inv_net;
    logic q_holder_net;

//////////////////////////////////////////////////////////////////////////////////////////////////
// COMBINATIONAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    assign clk_inv_net = ~clk_i;

    assign pll_o = q_holder_net & clk_i;

//////////////////////////////////////////////////////////////////////////////////////////////////
// SEQUENTIAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @ (posedge clk_inv_net or negedge arst_ni) begin
        if (~arst_ni) begin
            q_holder_net <= 0;
        end else begin
            q_holder_net <= en_i;
    end
    end



endmodule
