///////////////////////////////////////////////////////////////////////////////
//Author: Md Nazmus Sakib
//This is a delay generator which is constructed using counter
///////////////////////////////////////////////////////////////////////////////

module delay_gen #(
    parameter int COUNT_RANGE = 128
)(
    input  logic                  clk_i,
    input  logic                  arst_n_i,
    output logic                  delayed_o
);

//////////////////////////////////////////////////////////////////////////////////////////////////
// SIGNALS
//////////////////////////////////////////////////////////////////////////////////////////////////

    logic [$clog(n+1)-1:0] count_net;
    logic                  en_net;

//////////////////////////////////////////////////////////////////////////////////////////////////
// COMBINATIONAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    assign delayed_o=(count_net + 1 == COUNT_RANGE);
    assign en_net=~delayed_o;

//////////////////////////////////////////////////////////////////////////////////////////////////
// SEQUENTIAL
//////////////////////////////////////////////////////////////////////////////////////////////////

    always_ff @(posedge clk_i or negedge arst_n_i) begin
        if (arst_n_i) begin
            count_net <= 0;
        end else begin
            if(en) begin
                count_net <= count_net + 1;
            end
        end
    end

endmodule

